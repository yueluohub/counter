module counter_all ();
endmodule
