`timescale 1ns / 1ps 
module bfm_smartcard_iso7816(
    input wire i_clk;
    input wire i_rstn;
    inout wire io_data
);

parameter PARA_F=32'd372;
            PARA_D=32'd1;
            
















endmodule
